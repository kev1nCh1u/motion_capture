
module sources (
	probe);	

	input	[99:0]	probe;
endmodule
